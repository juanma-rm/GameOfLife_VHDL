----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- cells_tb.vhd
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
-- Import of libraries and packages
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.env.finish;

use work.utils_pkg.all;

----------------------------------------------------------------------------------
-- Entity
----------------------------------------------------------------------------------

entity cells_tb is
end;

----------------------------------------------------------------------------------
-- Architecture
----------------------------------------------------------------------------------

architecture bench of cells_tb is

    -- Constants


    -- Clock and reset

    constant clk_period_ns_c : time := 100 ns; -- 10 MHz
    signal clk_s    : std_ulogic := '0';
    signal rst_s    : std_ulogic := '0';

    -- dut signals

    signal   cells_arr_s : std_logic_vector(num_rows_c*num_cols_c - 1 downto 0);
    signal   done_s      : std_logic;
    signal   next_iter_s : std_logic;

begin

    --------------------------------------------------------------
    -- Clock and reset
    --------------------------------------------------------------

    clk_s <= not clk_s after clk_period_ns_c/2;
    rst_s <= '0', '1' after 10*clk_period_ns_c, '0' after 20*clk_period_ns_c;

    --------------------------------------------------------------
    -- Main process
    --------------------------------------------------------------

    process
    begin
        wait for 30 us;
        finish;                       
    end process;

    --------------------------------------------------------------
    -- DUT
    --------------------------------------------------------------

    cells_inst : entity work.cells
        port map (
            clk_i       => clk_s,
            rst_i       => rst_s,
            next_iter_i => next_iter_s,
            done_o      => done_s,
            cells_arr_o => cells_arr_s
        );
  
  
    --------------------------------------------------------------
    -- Stimulus
    --------------------------------------------------------------

    next_iter_s <= '1' when (done_s = '1') else '0';

    --------------------------------------------------------------
    -- Check
    --------------------------------------------------------------


end;
